-- ==============================================
--    Logic 3- to 8-Line Decoder/Demultiplexer
-- ==============================================
--
--                    CD74HC238
--                 +-------------+
--              3  |             |
--           >--/--|  A          |  8
--                 |          Y  |--/-->
--              3  |             |
--           >--/--| E           |
--                 |             |
--                 +-------------+
--
-- ===========
-- Truth table
-- ===========
--
-- See http://www.ti.com/lit/ds/symlink/cd74hc238.pdf
--
-- ==============================================

library ieee;
use ieee.std_logic_1164.all;

entity cd74hc238 is
    -- Declare interface based on the testbench spec.
end entity;

architecture behavioral of cd74hc238 is
begin
    -- Define behavioral architecture based on the CD74HC238 datasheet.
end architecture;
